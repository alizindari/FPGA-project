module instruction_mem #(parameter M=5, N=32) (input clk,
					       input [4:0] address,
					       output reg[31:0] instruction); 

reg [31:0] mem [0:31];


initial begin
//mem[0] =   32'b100000_00101_00000_0000000000000000;
mem[0] =   32'b111000_00000_00000_0000000000000111;
//mem[0] =   32'b110000_00000_00000_0000000000000111;
//mem[0] = 32'b001000_00000_00001_0000000000000011;
//mem[1] = 32'b001000_00000_00010_0000000000000011;
//mem[2] = 32'b000000_00001_00010_00011_00000_011000;
//mem[3] = 32'b100011_00010_00001_0000000000001010;
//mem[4] = 32'b000100_00001_00010_0000000000010100;
//mem[2] = 32'b000000_00001_00010_00011_00000_011000;
end

always @( posedge clk) begin 

	instruction <= mem[address];	
		
end 

endmodule
